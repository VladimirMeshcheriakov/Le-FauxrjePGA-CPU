// This file defines some opcodes of the ALU


`define AND   4'b0000
`define OR    4'b0001
`define ADD   4'b0010
`define XOR   4'b0011
`define SLL   4'b0100
`define SRL   4'b0101
`define SUB   4'b0110
`define SLT   4'b1001
`define SLTU  4'b1010
`define SLLI  4'b1100
`define SRLI  4'b1101
