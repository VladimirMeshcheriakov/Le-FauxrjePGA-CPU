// This file contains all the Store instruction definitons (the funct3 field)

`define SB 3'b000
`define SH 3'b001
`define SW 3'b010