// The cell_numbers parameter of the instruction_fetch.v is defined here:

`define CELL_NUMBERS   256