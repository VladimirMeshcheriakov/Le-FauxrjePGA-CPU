// This file defines some opcodes of the ALU


`define ADD   4'b0000
`define SLL    4'b0001
`define SLT   4'b0010
`define SLTU   4'b0011
`define XOR   4'b0100
`define SRL   4'b0101
`define OR   4'b0110
`define AND   4'b0111
`define SUB  4'b1000


