// This header file defines the branch operations

`define BEQ 3'b000
`define BNE 3'b001
`define JAL 3'b010
`define JALR 3'b011
`define BLT 3'b100
`define BGE 3'b101
`define BLTU 3'b110
`define BGEU 3'b111