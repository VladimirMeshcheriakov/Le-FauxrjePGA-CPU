// This file defines opcodes for the RISCV32I instruction types

`define U_TYPE_LUI      7'b0110111
`define U_TYPE_AUIPC    7'b0010111
`define J_TYPE_JAL      7'b1101111
`define I_TYPE_JALR     7'b1100111 
`define B_TYPE          7'b1100011
`define I_TYPE_LW       7'b0000011
`define S_TYPE          7'b0100011
`define I_TYPE_IMM      7'b0010011
`define R_TYPE          7'b0110011






